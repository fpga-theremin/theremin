.SUBCKT BB814/SIE 100 200 300
*anode1:         100
*anode2:         200
*common cathode: 300
*Package SOT23_2:
LIND1     1   10   0.77nH
LIND2     2   20   0.77nH
CAP2     10   20   73fF  
CAP3      3   10   120fF 
CAP4      3   20   120fF 
LIND10   10  100   0.56nH
LIND20   20  200   0.56nH
LIND30    3  300   0.49nH
*internal diodes:
D1 1 3 D1
D2 2 3 D1
R1 1 3 90e9
R2 2 3 90e9
.MODEL D1 D(IS=4.1f N=1.0 RS=260.0m XTI=3.5 EG=1.16
+ CJO=83.9p M=0.775 VJ=1.6 FC=0.5 TT=137.0n BV=33.5 IBV=1.0e-9)
.ENDS
