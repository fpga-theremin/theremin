.SUBCKT BB914 100 200 300
*anode1:         100
*anode2:         200
*common cathode: 300
*Package SOT23_2:
LIND1     1   10   0.77nH
LIND2     2   20   0.77nH
CAP2     10   20   73fF  
CAP3      3   10   120fF 
CAP4      3   20   120fF 
LIND10   10  100   0.56nH
LIND20   20  200   0.56nH
LIND30    3  300   0.49nH
*internal diodes:
D1 1 3 D1
D2 2 3 D1
R1 1 3 150e9
R2 2 3 150e9
.MODEL D1 D(IS=4.8f N=1.01 RS=280.0m XTI=3.0 EG=1.16
+ CJO=84.7873p M=0.819203 VJ=1.57986 FC=0.5 TT=137n BV=35.5 IBV=0.3e-9)
.ENDS
