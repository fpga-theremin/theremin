* AD8616 SPICE Macro-model
* Typical Values at Vs=�2.5V
* 05/04, Ver. 1.0
* Soufiane Bendaoud, ADSiV apps
*
* Copyright 2004 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of this
* model indicates your acceptance of the terms and provisions in
* the License Statement.
*
* Node Assignments
*			noninverting input
*			|	inverting input
*			|	|	 positive supply
*			|	|	 |	 negative supply
*			|	|	 |	 |	 output
*			|	|	 |	 |	 |
*			|	|	 |	 |	 |
.SUBCKT AD8616	1	2	99	50	45
* 
* INPUT STAGE
*
M1  14  7  8  8 PIX L=1E-6 W=1580E-6
M2  16  2  8  8 PIX L=1E-6 W=1580E-6
M3  17  7 10 10 NIX L=1E-6 W=1580E-6
M4  18  2 10 10 NIX L=1E-6 W=1580E-6
RC5 14 50 4E+3
RC6 16 50 4E+3
RC7 99 17 4E+3
RC8 99 18 4E+3
C1  14 16 0.08E-12
C2  17 18 0.08E-12
I1  99  8 100E-6
I2  10 50 100E-6
V1  99  9 0.2
V2  13 50 0.2
D1   8  9 DX
D2  13 10 DX
EOS  7  1 POLY(4) (22,98) (73,98) (81,98) (70,98) 23E-6 1 1 1 1
IOS  1  2  0.05E-12

*
*CMRR=100dB, ZERO AT 1MHz
*
 E1 21 98 POLY(2) (1,98) (2,98) 0 0.001255943   0.001255943
 R10 21 22 1.59E1
 R20 22 98 1.59E-1
 C10 21 22 1E-6

*
* PSRR=95dB, ZERO AT 534Hz
*
EPSY 98 72 POLY(1) (99,50) 0 0.5
CPS3 72 73 1E-6
RPS3 72 73 3.98E1
RPS4 73 98 7.96E-3
*
*
* VOLTAGE NOISE REFERENCE OF 8nV/rt(Hz)
*
VN1 80 98 0
RN1 80 98 16.45E-3
HN  81 98 VN1 7
RN2 81 98 1

*flicker noise 

D5 69 98 DNOISE
VSN 69 98 DC .6551
H1 70 98 VSN 25.3
RN 70 98 1

*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 .5 .5
GSY  99 50 (99,50) 240E-6 
EVP  97 98 POLY(1) (99,50) -0.6 0.5
EVN  51 98 POLY(1) (50,99) 0.6 0.5
*
* GAIN STAGE
*
G1 98 30 POLY(2) (14,16) (17,18) 0 2.1E-4 2.1E-4
R1 30 98 3.634E7
CF 45 30 14E-12
D3 30 97 DX
D4 51 30 DX
*
* OUTPUT STAGE
*
M5  45 46 99 99 POX L=1E-6 W=4.03E-3   
M6  45 47 50 50 NOX L=1E-6 W=4.03E-3  
EG1 99 46 POLY(1) (98,30) 0.45 1
EG2 47 50 POLY(1) (30,98) 0.45 1


*
* MODELS
*
.MODEL POX PMOS (LEVEL=2,KP=10E-6,VTO=-0.328,LAMBDA=0.01,RD=0)
.MODEL NOX NMOS (LEVEL=2,KP=10E-6,VTO=+0.328,LAMBDA=0.01,RD=0)
.MODEL PIX PMOS (LEVEL=2,KP=10E-6,VTO=-0.328,LAMBDA=0.01,TOX=100E-3)
.MODEL NIX NMOS (LEVEL=2,KP=10E-6,VTO=+0.328,LAMBDA=0.01,TOX=100E-3)
.MODEL DX D(IS=1E-14,RS=5,KF=1E-15)
.MODEL DNOISE D(IS=1E-14,RS=0,KF=1E-15)

.ENDS AD8616
*
*$

*$
