module theremin_io_ip_tb();


endmodule;
