* ADG721 SPICE Macro-model
* Generic Desc:CMOS, Low Voltage, 4 Ohm Dual SPST Switches in 3 mm x 2 mm LFCSP
* Developed by: mbarrien / ANALOG
* Revision History: 2.0 (8/2018) - Updated model design
* 1.2 (05/2008)
* Copyright 2018 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement. Use of this model 
* indicates your acceptance of the terms and provisions in the License Statement.
*
* Begin Notes:
* The model will work on Vdd from 0.5V to 5V single supply.
* The model provides parametric specifications at 5V only and is not variable with Vdd changes. Please see datasheet spec table.
*
* Parameters modeled include:
* On Resistance
* Ton and Toff
* Break-Before-Make
* Off Isolation
* Crosstalk
* Supply Currents: Iss/Idd
* Bandwidth
* Charge Injection
* Connections
*      1  = S1
*      2  = D1
*      3  = IN2
*      4  = GND
*      5  = S2
*      6  = D2
*      7  = IN1
*      8  = VDD
*
.SUBCKT ADG721 1 2 3 4 5 6 7 8

.MODEL VON VSWITCH(Von=5 Voff=0.8 Ron=0.001 Roff=9000000000000)
.MODEL VEN VSWITCH(Von=5 Voff=0.8 Ron=7100 Roff=23000)
.MODEL VRESET VSWITCH(Von=5 Voff=0.8 Ron=2700000 Roff=1000)
.MODEL DCLAMP D(IS=1E-15 IBV=1E-13)


* CROSSTALK
C12X 1 5 44E-015

* IDD/ISS
I1 8 4 0.001E-006

* Configuration: SPST 2:2


** SWITCH 1 **
*
* ESD PROTECTION DIODES
D11 4 2 DCLAMP
D12 2 8 DCLAMP
D13 4 1 DCLAMP
D14 1 8 DCLAMP
*
* OFF ISOLATION
C11 1 2 0.32E-012
*
* CHARGE INJECTION
C12 2 140 0.62E-012
C13 1 140 0.62E-012
*
* CD/CS OFF AND BANDWIDTH
C14 1 4 12.75E-012
C15 2 4 12.75E-012
*
* ON RESISTANCE
Ech155 1555 4 VALUE = { IF ((ABS(V(1)))>(ABS(V(184))),V(1),V(2)) }
R155 1555 4 1G
R11 137 2 0.001
S111 136 141 1141 4 VON
Ech111 1141 4 VALUE = { IF (V(1555)<1.2,5,0) }
Ech11 141 4 VALUE = { IF (V(1555)<1.2,0.291666666666667*(V(1555)-1.2)+3.15,0) }
S112 136 146 1146 4 VON
Ech112 1146 4 VALUE = { IF ((V(1555)>=1.2) & (V(1555)<=3.75),5,0) }
Ech12 146 4 VALUE = { IF ((V(1555)>=1.2) & (V(1555)<=3.75),((3.15-2.8)/((1.2-2.30422720885496)*(1.2-2.30422720885496)))*(V(1555)-2.30422720885496)*(V(1555)-2.30422720885496) + 2.8,0) }
S113 136 144 1144 4 VON
Ech113 1144 4 VALUE = { IF (V(1555)>3.75,5,0) }
Ech13 144 4 VALUE = { IF (V(1555)>3.75,-0.264*(V(1555)-3.75)+3.4,0) }
RIN1	136 4	1G
EOUT1 137 181	POLY(2) (136,4) (180,4) 0 0 0 0 0.999/1000
FCOPY1	4 180 VSENSE1 1
RSENSOR1 180 4	1K
VSENSE1 181 184	0
*
* TON/ TOFF/ BBM
S11 182 184 140 4 VON
S12 143 138 143 4 VEN
Ech14 143 4 VALUE = { IF(V(7)>=2.4, 5 , 0.8 ) }
eV1 140 4 138 4 1
C16 138 4 1e-012
*
* VOLTAGE SUPPLY REQUIREMENT
S13 1 182 185 4 VON
S15 139 185 139 4 VON
Ech16 139 4 VALUE = { IF((V(0)>=-0.5 & (V(8)<=5 & V(8)>=0.5)), 5 , 0.01 ) }


** SWITCH 2 **
*
* ESD PROTECTION DIODES
D21 0 6 DCLAMP
D22 6 8 DCLAMP
D23 0 5 DCLAMP
D24 5 8 DCLAMP
*
* OFF ISOLATION
C21 5 6 0.32E-012
*
* CHARGE INJECTION
C22 6 240 0.62E-012
C23 5 240 0.62E-012
*
* CD/CS OFF AND BANDWIDTH
C24 5 4 12.75E-012
C25 6 4 12.75E-012
*
* ON RESISTANCE
Ech255 2555 4 VALUE = { IF ((ABS(V(5)))>(ABS(V(284))),V(5),V(6)) }
R255 2555 4 1G
R21 237 6 0.001
S221 236 241 2241 4 VON
Ech221 2241 4 VALUE = { IF (V(2555)<1.2,5,0) }
Ech21 241 4 VALUE = { IF (V(2555)<1.2,0.291666666666667*(V(2555)-1.2)+3.15,0) }
S222 236 246 2246 4 VON
Ech222 2246 4 VALUE = { IF ((V(2555)>=1.2) & (V(2555)<=3.75),5,0) }
Ech22 246 4 VALUE = { IF ((V(2555)>=1.2) & (V(2555)<=3.75),((3.15-2.8)/((1.2-2.30422720885496)*(1.2-2.30422720885496)))*(V(2555)-2.30422720885496)*(V(2555)-2.30422720885496) + 2.8,0) }
S223 236 244 2244 4 VON
Ech223 2244 4 VALUE = { IF (V(2555)>3.75,5,0) }
Ech23 244 4 VALUE = { IF (V(2555)>3.75,-0.264*(V(2555)-3.75)+3.4,0) }
RIN2	236 4	1G
EOUT2 237 281	POLY(2) (236,4) (280,4) 0 0 0 0 0.999/1000
FCOPY2	4 280 VSENSE2 1
RSENSOR2 280 4	1K
VSENSE2 281 284	0
*
* TON/ TOFF/ BBM
S21 282 284 240 4 VON
S22 243 238 243 4 VEN
Ech24 243 4 VALUE = { IF(V(3)>=2.4, 5 , 0.8 ) }
eV2 240 4 238 4 1
C26 238 4 1e-012
*
* VOLTAGE SUPPLY REQUIREMENT
S23 5 282 285 4 VON
S25 239 285 239 4 VON
Ech26 239 4 VALUE = { IF((V(0)>=-0.5 & (V(8)<=5 & V(8)>=0.5)), 5 , 0.01 ) }

.ENDS ADG721
